`define NUM_STATES 256 

module microstore(output reg[39:0] out,
                  output reg [9:0] current_state,
                  input[9:0] next_state,
                  input reset);
/* state_info contains control signal bits for all states. **state_info[0] corresponds to State 0, state_info[1] to State 1, etc.**
 **MUST FILL UNUSED STATES WITH ZEROS SO ARRAY POSITIONS CORRESPOND TO THEIR STATE***/
parameter[0:40 * `NUM_STATES - 1] state_info = {
40'h2100334c00,
40'h6040813c00,
40'h611c835800,
40'hb09c000003,
40'h9400000001,
40'h0000000000, // 5
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h2300100000,
40'h2100100000,
40'h2100930000,
40'h4100873c0c,
40'h0000000000, 
40'h0000000000, // 15
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h4040118028,
40'h4040018028,
40'h4140158028,
40'h4140058028,
40'h604001bc00,
40'h602041bc00,
40'h410815802a,
40'h604001bc00,
40'h602041bc00,
40'h410805802a,
40'h4040118828,
40'h4040018828,
40'h4140158828,
40'h4140058828,
40'h604001bc00,
40'h602041bc00,
40'h410815882a,
40'h604001bc00,
40'h602041bc00,
40'h410805882a,
40'h602041bc00,
40'h6008018000,
40'hf00801802a,
40'h404411803f,
40'h404401803f,
40'h414415803f,
40'h414405803f,
40'h604401bc00,
40'h602441bc00,
40'h410c158041,
40'h604401bc00,
40'h602441bc00,
40'h410c058041,
40'h404411883f,
40'h404401883f,
40'h414415883f,
40'h414405883f,
40'h604401bc00,
40'h602441bc00,
40'h410c158841,
40'h604401bc00,
40'h602441bc00,
40'h410c058841,
40'h602441bc00,
40'h600c018000,
40'hf00c018041,
40'h4040110052,
40'h4040010052,
40'h4140150052,
40'h4140050052,
40'h6040013c00,
40'h4100150052,
40'h6040013c00,
40'h4100050052,
40'h4040110852,
40'h4040010852,
40'h4140150852,
40'h4140050852,
40'h6040013c00,
40'h4100150852,
40'h6040013c00,
40'h4100050852,
40'h6018010000,
40'hb038010053,
40'h2100214c00,
40'h4044110065,
40'h4044010065,
40'h4144150065,
40'h4144050065,
40'h6044013c00,
40'h4104150065,
40'h6044013c00,
40'h4104050065,
40'h4044110865,
40'h4044010865,
40'h4144150865,
40'h4144050865,
40'h6044013c00,
40'h4104150865,
40'h6044013c00,
40'h4104050865,
40'h601c010000,
40'hb03c010066,
40'h2104214c00,
40'h404211807c,
40'h404201807c,
40'h414215807c,
40'h414205807c,
40'h604201bc00,
40'h602241bc00,
40'h410a15807e,
40'h604201bc00,
40'h602241bc00,
40'h410a05807c,
40'h404211887c,
40'h404201887c,
40'h414215887c,
40'h414205887c,
40'h604201bc00,
40'h602241bc00,
40'h410a15887e,
40'h604201bc00,
40'h602241bc00,
40'h410a05887e,
40'h602241bc00,
40'h600a018000,
40'hf00a01807e,
40'h404211008f,
40'h404201008f,
40'h414215008f,
40'h414205008f,
40'h6042013c00,
40'h410215008f,
40'h6042013c00,
40'h410205008f,
40'h404211088f,
40'h404201088f,
40'h414215088f,
40'h414205088f,
40'h6042013c00,
40'h410215088f,
40'h6042013c00,
40'h410205088f,
40'h601a010000,
40'hb03a010090,
40'h2102214c00,
40'h40411100a2,
40'h40410100a2,
40'h41411500a2,
40'h41410500a2,
40'h6041013c00,
40'h41011500a2,
40'h6041013c00,
40'h41010500a2,
40'h40411108a2,
40'h40410108a2,
40'h41411508a2,
40'h41410508a2,
40'h6041013c00,
40'h41011508a2,
40'h6041013c00,
40'h41010508a2,
40'h6019010000,
40'hb0390100a3,
40'h2101214c00,
40'h40431100b5,
40'h40430100b5,
40'h41431500b5,
40'h41430500b5,
40'h6043013c00,
40'h41031500b5,
40'h6043013c00,
40'h41030500b5,
40'h40431108b5,
40'h40430108b5,
40'h41431508b5,
40'h41430508b5,
40'h6043013c00,
40'h41031508b5,
40'h6043013c00,
40'h41030508b5,
40'h601b010000,
40'hb03b0100b6,
40'h2103214c00,
40'h40441100c8,
40'h40440100c8,
40'h41441500c8,
40'h41440500c8,
40'h6044013c00,
40'h41041500c8,
40'h6044013c00,
40'h41040500c8,
40'h40441108c8,
40'h40440108c8,
40'h41441508c8,
40'h41440508c8,
40'h6044013c00,
40'h41041508c8,
40'h6044013c00,
40'h41040508c8,
40'h601c010000,
40'hb03c0100c9,
40'h6104214c00,
40'h6044115c00,
40'h601c010000,
40'hb03c0100cd,
40'h2104294c00,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000
};

integer i;

always @(next_state, reset)
begin
    if (reset) begin
        out           <= state_info[0+:40];
        current_state <= 10'd0;
    end
    else begin
        out           <= state_info[40*next_state+:40];
        current_state <= next_state;
    end
end

endmodule
