module binary_decoder_test;

endmodule