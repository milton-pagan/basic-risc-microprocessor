module shift_sign_extender_test();
    
    wire[31:0] out;
    wire carry_out;
    
    reg[31:0] instruction, Rm;
    
endmodule
