module conditions_mux(output reg out,
                      input in0,
                      in1,
                      in2,
                      in3,
                      input[1:0] select);

                      
    
endmodule
