`define NUM_STATES 256 

module microstore(output reg[38:0] out,
                  output reg [9:0] current_state,
                  input[9:0] next_state,
                  input reset);
/* state_info contains control signal bits for all states. **state_info[0] corresponds to State 0, state_info[1] to State 1, etc.**
 **MUST FILL UNUSED STATES WITH ZEROS SO ARRAY POSITIONS CORRESPOND TO THEIR STATE***/
parameter[0:39 * `NUM_STATES - 1] state_info = {
39'h10801b4c00, // 0
39'h3020413c00,
39'h308e435800,
39'h584e000003,
39'h4a00000001,
39'h0000000000, // 5
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h1180080000, // 10
39'h1080080000,
39'h10804b5c00,
39'h2080473c0c,
39'h0000000000, 
39'h0000000000, // 15
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h2020098028, // 20
39'h2020018028,
39'h20a00d8028,
39'h20a0058028,
39'h302001bc00,
39'h301021bc00, // 25
39'h20840d802a,
39'h302001bc00,
39'h301021bc00,
39'h208405802a,
39'h2020098828, // 30
39'h2020018828,
39'h20a00d8828,
39'h20a0058828,
39'h302001bc00,
39'h301021bc00, // 35
39'h20840d882a,
39'h302001bc00,
39'h301021bc00,
39'h208405882a,
39'h301021bc00, // 40
39'h3004018000,
39'h780401802a,
39'h202209803f,
39'h202201803f,
39'h20a20d803f, // 45
39'h20a205803f,
39'h302201bc00,
39'h301221bc00,
39'h20860d8041,
39'h302201bc00, // 50
39'h301221bc00,
39'h2086058041,
39'h202209883f,
39'h202201883f,
39'h20a20d883f, // 55
39'h20a205883f,
39'h302201bc00,
39'h301221bc00,
39'h20860d8841,
39'h302201bc00, // 60
39'h301221bc00,
39'h2086058841,
39'h301221bc00,
39'h3006018000,
39'h7806018041, // 65
39'h2020090052,
39'h2020010052,
39'h20a00d0052,
39'h20a0050052,
39'h3020013c00, // 70
39'h20800d0052,
39'h3020013c00,
39'h2080050052,
39'h2020090852,
39'h2020010852, // 75
39'h20a00d0852,
39'h20a0050852,
39'h3020013c00,
39'h20800d0852,
39'h3020013c00, // 80
39'h2080050852,
39'h300c010000,
39'h581c010053,
39'h1080114c00,
39'h2022090065, // 85
39'h2022010065,
39'h20a20d0065,
39'h20a2050065,
39'h3022013c00,
39'h20820d0065, // 90
39'h3022013c00,
39'h2082050065,
39'h2022090865,
39'h2022010865,
39'h20a20d0865, // 95
39'h20a2050865,
39'h3022013c00,
39'h20820d0865,
39'h3022013c00,
39'h2082050865, // 110
39'h300e010000,
39'h581e010066,
39'h1082114c00,
39'h202189807c,
39'h202181807c, // 105
39'h20a18d807c,
39'h20a185807c,
39'h302181bc00,
39'h3011a1bc00,
39'h20858d807e, // 110
39'h302181bc00,
39'h3011a1bc00,
39'h208585807c,
39'h202189887c,
39'h202181887c, // 115
39'h20a18d887c,
39'h20a185887c,
39'h302181bc00,
39'h3011a1bc00,
39'h20858d887e, // 120
39'h302181bc00,
39'h3011a1bc00,
39'h208585887e,
39'h3011a1bc00,
39'h3005818000, // 125
39'h780581807e,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000,
39'h0000000000
};

integer i;

always @(next_state, reset)
begin
    if (reset) begin
        out           <= state_info[0+:39];
        current_state <= 10'd0;
    end
    else begin
        out           <= state_info[39*next_state+:39];
        current_state <= next_state;
    end
end

endmodule
