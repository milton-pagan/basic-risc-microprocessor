`define NUM_STATES 256 

module microstore(output reg[39:0] out,
                  output reg [9:0] current_state,
                  input[9:0] next_state,
                  input reset);
/* state_info contains control signal bits for all states. **state_info[0] corresponds to State 0, state_info[1] to State 1, etc.**
 **MUST FILL UNUSED STATES WITH ZEROS SO ARRAY POSITIONS CORRESPOND TO THEIR STATE***/
parameter[0:40 * `NUM_STATES - 1] state_info = {
40'h2100333400,
40'h6040814000,
40'h611c834400,
40'hb09c001003,
40'h9400001001,
40'h0000000000, // 5
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h2300101000,
40'h2100101000,
40'h2100931000,
40'h410087400c,
40'h2200101000,
40'h0000000000, // 15
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h4040119028,
40'h4040019028,
40'h4140159028,
40'h4140059028,
40'h604001c000,
40'h602041c000,
40'h410815902a,
40'h604001c000,
40'h602041c000,
40'h410805902a,
40'h4040118828,
40'h4040018828,
40'h4140158828,
40'h4140058828,
40'h604001c000,
40'h602041c000,
40'h410815882a,
40'h604001c000,
40'h602041c000,
40'h410805882a,
40'h602041c000,
40'h6008019000,
40'hf00801902a,
40'h404411903f,
40'h404401903f,
40'h414415903f,
40'h414405903f,
40'h604401c000,
40'h602441c000,
40'h410c159041,
40'h604401c000,
40'h602441c000,
40'h410c059041,
40'h404411883f,
40'h404401883f,
40'h414415883f,
40'h414405883f,
40'h604401c000,
40'h602441c000,
40'h410c158841,
40'h604401c000,
40'h602441c000,
40'h410c058841,
40'h602441c000,
40'h600c019000,
40'hf00c019041,
40'h4040111052,
40'h4040011052,
40'h4140151052,
40'h4140051052,
40'h6040014000,
40'h4100151052,
40'h6040014000,
40'h4100050052,
40'h4040110852,
40'h4040010852,
40'h4140150852,
40'h4140050852,
40'h6040014000,
40'h4100150852,
40'h6040014000,
40'h4100050852,
40'h6018011000,
40'hb038011053,
40'h2100213400,
40'h4044111065,
40'h4044011065,
40'h4144151065,
40'h4144051065,
40'h6044014000,
40'h4104151065,
40'h6044014000,
40'h4104051065,
40'h4044110865,
40'h4044010865,
40'h4144150865,
40'h4144050865,
40'h6044014000,
40'h4104150865,
40'h6044014000,
40'h4104050865,
40'h601c011000,
40'hb03c011066,
40'h2104213400,
40'h404211907c,
40'h404201907c,
40'h414215907c,
40'h414205907c,
40'h604201c000,
40'h602241c000,
40'h410a15907e,
40'h604201c000,
40'h602241c000,
40'h410a05907c,
40'h404211887c,
40'h404201887c,
40'h414215887c,
40'h414205887c,
40'h604201c000,
40'h602241c000,
40'h410a15887e,
40'h604201c000,
40'h602241c000,
40'h410a05887e,
40'h602241c000,
40'h600a019000,
40'hf00a01907e,
40'h404211108f,
40'h404201108f,
40'h414215108f,
40'h414205108f,
40'h6042014000,
40'h410215108f,
40'h6042014000,
40'h410205108f,
40'h404211088f,
40'h404201088f,
40'h414215088f,
40'h414205088f,
40'h6042014000,
40'h410215088f,
40'h6042014000,
40'h410205088f,
40'h601a011000,
40'hb03a011090,
40'h2102213400,
40'h40411110a2,
40'h40410110a2,
40'h41411510a2,
40'h41410510a2,
40'h6041014000,
40'h41011510a2,
40'h6041014000,
40'h41010510a2,
40'h40411108a2,
40'h40410108a2,
40'h41411508a2,
40'h41410508a2,
40'h6041014000,
40'h41011508a2,
40'h6041014000,
40'h41010508a2,
40'h6019011000,
40'hb0390110a3,
40'h2101213400,
40'h40431110b5,
40'h40430110b5,
40'h41431510b5,
40'h41430510b5,
40'h6043014000,
40'h41031510b5,
40'h6043014000,
40'h41030510b5,
40'h40431108b5,
40'h40430108b5,
40'h41431508b5,
40'h41430508b5,
40'h6043014000,
40'h41031508b5,
40'h6043014000,
40'h41030508b5,
40'h601b011000,
40'hb03b0110b6,
40'h2103213400,
40'h40441110c8,
40'h40440110c8,
40'h41441510c8,
40'h41440510c8,
40'h6044014000,
40'h41041510c8,
40'h6044014000,
40'h41040510c8,
40'h40441108c8,
40'h40440108c8,
40'h41441508c8,
40'h41440508c8,
40'h6044014000,
40'h41041508c8,
40'h6044014000,
40'h41040508c8,
40'h601c011000,
40'hb03c0110c9,
40'h6104213400,
40'h6044114800,
40'h601c011000,
40'hb03c0110cd,
40'h2104293400,
40'h40441190e3,
40'h40440190e3,
40'h41441590e3,
40'h41440590e3,
40'h604401c000,
40'h602441c000,
40'h410c1590e5,
40'h604401c000,
40'h602441c000,
40'h410c0590e5,
40'h40441188e3,
40'h40440188e3,
40'h41441588e3,
40'h41440588e3,
40'h604401c000,
40'h602441c000,
40'h410c1588e5,
40'h604401c000,
40'h602441c000,
40'h410c0588e5,
40'h602441c000,
40'h600c019000,
40'hb00c0190e5,
40'h604411c800,
40'h6024c1c000,
40'h600c019000,
40'hf00c0190e9,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000,
40'h0000000000
};

integer i;

always @(next_state, reset)
begin
    if (reset) begin
        out           <= state_info[0+:40];
        current_state <= 10'd0;
    end
    else begin
        out           <= state_info[40*next_state+:40];
        current_state <= next_state;
    end
end

endmodule
